`timescale 1ns / 1ps

module prop(output p ,input a, b);
    assign p=a^b;
endmodule
