`timescale 1ns / 1ps
module gen(output  g,input  a,b);
   assign g=a&b;   
endmodule